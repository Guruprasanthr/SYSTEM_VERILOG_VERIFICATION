interface intf;
  logic clk;
  logic rst;
  logic up;
  logic [3:0]count;
endinterface
  
